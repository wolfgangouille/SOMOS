`timescale 1ns / 1ps

module COVAR_8(M_CLK,TRIGGER,NEW_DATA1,NEW_DATA2,NEW_DATA3,NEW_DATA4,NEW_DATA5,NEW_DATA6,NEW_DATA7,NEW_DATA8,COVAR11,COVAR22,COVAR33,COVAR44,COVAR55,COVAR66,COVAR77,COVAR88,DATA_READY);

input TRIGGER;
input [15:0] NEW_DATA1;
input [15:0] NEW_DATA2;
input [15:0] NEW_DATA3;
input [15:0] NEW_DATA4;
input [15:0] NEW_DATA5;
input [15:0] NEW_DATA6;
input [15:0] NEW_DATA7;
input [15:0] NEW_DATA8;
input M_CLK;

output [15:0] COVAR11;
output [15:0] COVAR22;
output [15:0] COVAR33;
output [15:0] COVAR44;
output [15:0] COVAR55;
output [15:0] COVAR66;
output [15:0] COVAR77;
output [15:0] COVAR88;

/*output [15:0] COVAR12;
output [15:0] COVAR13;
output [15:0] COVAR14;
output [15:0] COVAR15;
output [15:0] COVAR16;
output [15:0] COVAR17;
output [15:0] COVAR18;
output [15:0] COVAR23;
output [15:0] COVAR24;
output [15:0] COVAR25;
output [15:0] COVAR26;
output [15:0] COVAR27;
output [15:0] COVAR28;
output [15:0] COVAR34;
output [15:0] COVAR35;
output [15:0] COVAR36;
output [15:0] COVAR37;
output [15:0] COVAR38;
output [15:0] COVAR45;
output [15:0] COVAR46;
output [15:0] COVAR47;
output [15:0] COVAR48;
output [15:0] COVAR56;
output [15:0] COVAR57;
output [15:0] COVAR58;
output [15:0] COVAR67;
output [15:0] COVAR68;
output [15:0] COVAR78;*/

output DATA_READY;

reg [15:0] DATA1;
reg [15:0] DATA2;
reg [15:0] DATA3;
reg [15:0] DATA4;
reg [15:0] DATA5;
reg [15:0] DATA6;
reg [15:0] DATA7;
reg [15:0] DATA8;

reg [31:0] TEMP_MEAN1;
reg [31:0] TEMP_MEAN2;
reg [31:0] TEMP_MEAN3;
reg [31:0] TEMP_MEAN4;
reg [31:0] TEMP_MEAN5;
reg [31:0] TEMP_MEAN6;
reg [31:0] TEMP_MEAN7;
reg [31:0] TEMP_MEAN8;

reg [15:0] MEAN1;
reg [15:0] MEAN2;
reg [15:0] MEAN3;
reg [15:0] MEAN4;
reg [15:0] MEAN5;
reg [15:0] MEAN6;
reg [15:0] MEAN7;
reg [15:0] MEAN8;

reg [15:0] DELTA_ABS1;
reg [15:0] DELTA_ABS2;
reg [15:0] DELTA_ABS3;
reg [15:0] DELTA_ABS4;
reg [15:0] DELTA_ABS5;
reg [15:0] DELTA_ABS6;
reg [15:0] DELTA_ABS7;
reg [15:0] DELTA_ABS8;

reg  DELTA_1_NEG;
reg  DELTA_2_NEG;
reg  DELTA_3_NEG;
reg  DELTA_4_NEG;
reg  DELTA_5_NEG;
reg  DELTA_6_NEG;
reg  DELTA_7_NEG;
reg  DELTA_8_NEG;

//Instantaneous covar??
reg [31:0] S11;
reg [31:0] S12;
reg [31:0] S13;
reg [31:0] S14;
reg [31:0] S15;
reg [31:0] S16;
reg [31:0] S17;
reg [31:0] S18;
reg [31:0] S22;
reg [31:0] S23;
reg [31:0] S24;
reg [31:0] S25;
reg [31:0] S26;
reg [31:0] S27;
reg [31:0] S28;
reg [31:0] S33;
reg [31:0] S34;
reg [31:0] S35;
reg [31:0] S36;
reg [31:0] S37;
reg [31:0] S38;
reg [31:0] S44;
reg [31:0] S45;
reg [31:0] S46;
reg [31:0] S47;
reg [31:0] S48;
reg [31:0] S55;
reg [31:0] S56;
reg [31:0] S57;
reg [31:0] S58;
reg [31:0] S66;
reg [31:0] S67;
reg [31:0] S68;
reg [31:0] S77;
reg [31:0] S78;
reg [31:0] S88;

reg [15:0] COVAR11;
reg [15:0] COVAR12;
reg [15:0] COVAR13;
reg [15:0] COVAR14;
reg [15:0] COVAR15;
reg [15:0] COVAR16;
reg [15:0] COVAR17;
reg [15:0] COVAR18;
reg [15:0] COVAR22;
reg [15:0] COVAR23;
reg [15:0] COVAR24;
reg [15:0] COVAR25;
reg [15:0] COVAR26;
reg [15:0] COVAR27;
reg [15:0] COVAR28;
reg [15:0] COVAR33;
reg [15:0] COVAR34;
reg [15:0] COVAR35;
reg [15:0] COVAR36;
reg [15:0] COVAR37;
reg [15:0] COVAR38;
reg [15:0] COVAR44;
reg [15:0] COVAR45;
reg [15:0] COVAR46;
reg [15:0] COVAR47;
reg [15:0] COVAR48;
reg [15:0] COVAR55;
reg [15:0] COVAR56;
reg [15:0] COVAR57;
reg [15:0] COVAR58;
reg [15:0] COVAR66;
reg [15:0] COVAR67;
reg [15:0] COVAR68;
reg [15:0] COVAR77;
reg [15:0] COVAR78;
reg [15:0] COVAR88;

reg [31:0] TEMP_COVAR11;
reg [31:0] TEMP_COVAR12;
reg [31:0] TEMP_COVAR13;
reg [31:0] TEMP_COVAR14;
reg [31:0] TEMP_COVAR15;
reg [31:0] TEMP_COVAR16;
reg [31:0] TEMP_COVAR17;
reg [31:0] TEMP_COVAR18;
reg [31:0] TEMP_COVAR22;
reg [31:0] TEMP_COVAR23;
reg [31:0] TEMP_COVAR24;
reg [31:0] TEMP_COVAR25;
reg [31:0] TEMP_COVAR26;
reg [31:0] TEMP_COVAR27;
reg [31:0] TEMP_COVAR28;
reg [31:0] TEMP_COVAR33;
reg [31:0] TEMP_COVAR34;
reg [31:0] TEMP_COVAR35;
reg [31:0] TEMP_COVAR36;
reg [31:0] TEMP_COVAR37;
reg [31:0] TEMP_COVAR38;
reg [31:0] TEMP_COVAR44;
reg [31:0] TEMP_COVAR45;
reg [31:0] TEMP_COVAR46;
reg [31:0] TEMP_COVAR47;
reg [31:0] TEMP_COVAR48;
reg [31:0] TEMP_COVAR55;
reg [31:0] TEMP_COVAR56;
reg [31:0] TEMP_COVAR57;
reg [31:0] TEMP_COVAR58;
reg [31:0] TEMP_COVAR66;
reg [31:0] TEMP_COVAR67;
reg [31:0] TEMP_COVAR68;
reg [31:0] TEMP_COVAR77;
reg [31:0] TEMP_COVAR78;
reg [31:0] TEMP_COVAR88;


reg [15:0] ALPHA_MEAN;
reg [15:0] ALPHA_RMS;

reg [1:0] TRIGSHIFT;
reg DATA_READY;

reg [7:0] COUNTER;

initial begin
	ALPHA_MEAN<=16'b0000000000000001;
	ALPHA_RMS<=16'b0000000000000100;

	DATA1<=16'b0;
	DATA2<=16'b0;
	DATA3<=16'b0;
	DATA4<=16'b0;
	DATA5<=16'b0;
	DATA6<=16'b0;
	DATA7<=16'b0;
	DATA8<=16'b0;

	TEMP_MEAN1<=32'b10000000000000000000000000000000;
	TEMP_MEAN2<=32'b10000000000000000000000000000000;
	TEMP_MEAN3<=32'b10000000000000000000000000000000;
	TEMP_MEAN4<=32'b10000000000000000000000000000000;
	TEMP_MEAN5<=32'b10000000000000000000000000000000;
	TEMP_MEAN6<=32'b10000000000000000000000000000000;
	TEMP_MEAN7<=32'b10000000000000000000000000000000;
	TEMP_MEAN8<=32'b10000000000000000000000000000000;



	MEAN1<=16'b0000000000000000;
	MEAN2<=16'b0000000000000000;
	MEAN3<=16'b0000000000000000;
	MEAN4<=16'b0000000000000000;
	MEAN5<=16'b0000000000000000;
	MEAN6<=16'b0000000000000000;
	MEAN7<=16'b0000000000000000;
	MEAN8<=16'b0000000000000000;


	DELTA_ABS1<=16'b0;
	DELTA_ABS2<=16'b0;
	DELTA_ABS3<=16'b0;
	DELTA_ABS4<=16'b0;
	DELTA_ABS5<=16'b0;
	DELTA_ABS6<=16'b0;
	DELTA_ABS7<=16'b0;
	DELTA_ABS8<=16'b0;

	DELTA_1_NEG<=1'b0;
	DELTA_2_NEG<=1'b0;
	DELTA_3_NEG<=1'b0;
	DELTA_4_NEG<=1'b0;
	DELTA_5_NEG<=1'b0;
	DELTA_6_NEG<=1'b0;
	DELTA_7_NEG<=1'b0;
	DELTA_8_NEG<=1'b0;


	S11<=32'b0;
	S12<=32'b0;
	S13<=32'b0;
	S14<=32'b0;
	S15<=32'b0;
	S16<=32'b0;
	S17<=32'b0;
	S18<=32'b0;
	S22<=32'b0;
	S23<=32'b0;
	S24<=32'b0;
	S25<=32'b0;
	S26<=32'b0;
	S27<=32'b0;
	S28<=32'b0;
	S33<=32'b0;
	S34<=32'b0;
	S35<=32'b0;
	S36<=32'b0;
	S37<=32'b0;
	S38<=32'b0;
	S44<=32'b0;
	S45<=32'b0;
	S46<=32'b0;
	S47<=32'b0;
	S48<=32'b0;
	S55<=32'b0;
	S56<=32'b0;
	S57<=32'b0;
	S58<=32'b0;
	S66<=32'b0;
	S67<=32'b0;
	S68<=32'b0;
	S77<=32'b0;
	S78<=32'b0;
	S88<=32'b0;


	COVAR11<=16'b0000000000000000;
	COVAR12<=16'b0000000000000000;
	COVAR13<=16'b0000000000000000;
	COVAR14<=16'b0000000000000000;
	COVAR15<=16'b0000000000000000;
	COVAR16<=16'b0000000000000000;
	COVAR17<=16'b0000000000000000;
	COVAR18<=16'b0000000000000000;
	COVAR22<=16'b0000000000000000;
	COVAR23<=16'b0000000000000000;
	COVAR24<=16'b0000000000000000;
	COVAR25<=16'b0000000000000000;
	COVAR26<=16'b0000000000000000;
	COVAR27<=16'b0000000000000000;
	COVAR28<=16'b0000000000000000;
	COVAR33<=16'b0000000000000000;
	COVAR34<=16'b0000000000000000;
	COVAR35<=16'b0000000000000000;
	COVAR36<=16'b0000000000000000;
	COVAR37<=16'b0000000000000000;
	COVAR38<=16'b0000000000000000;
	COVAR44<=16'b0000000000000000;
	COVAR45<=16'b0000000000000000;
	COVAR46<=16'b0000000000000000;
	COVAR47<=16'b0000000000000000;
	COVAR48<=16'b0000000000000000;
	COVAR55<=16'b0000000000000000;
	COVAR56<=16'b0000000000000000;
	COVAR57<=16'b0000000000000000;
	COVAR58<=16'b0000000000000000;
	COVAR66<=16'b0000000000000000;
	COVAR67<=16'b0000000000000000;
	COVAR68<=16'b0000000000000000;
	COVAR77<=16'b0000000000000000;
	COVAR78<=16'b0000000000000000;
	COVAR88<=16'b0000000000000000;



	TEMP_COVAR11<=32'b0;
	TEMP_COVAR12<=32'b0;
	TEMP_COVAR13<=32'b0;
	TEMP_COVAR14<=32'b0;
	TEMP_COVAR15<=32'b0;
	TEMP_COVAR16<=32'b0;
	TEMP_COVAR17<=32'b0;
	TEMP_COVAR18<=32'b0;
	TEMP_COVAR22<=32'b0;
	TEMP_COVAR23<=32'b0;
	TEMP_COVAR24<=32'b0;
	TEMP_COVAR25<=32'b0;
	TEMP_COVAR26<=32'b0;
	TEMP_COVAR27<=32'b0;
	TEMP_COVAR28<=32'b0;
	TEMP_COVAR33<=32'b0;
	TEMP_COVAR34<=32'b0;
	TEMP_COVAR35<=32'b0;
	TEMP_COVAR36<=32'b0;
	TEMP_COVAR37<=32'b0;
	TEMP_COVAR38<=32'b0;
	TEMP_COVAR44<=32'b0;
	TEMP_COVAR45<=32'b0;
	TEMP_COVAR46<=32'b0;
	TEMP_COVAR47<=32'b0;
	TEMP_COVAR48<=32'b0;
	TEMP_COVAR55<=32'b0;
	TEMP_COVAR56<=32'b0;
	TEMP_COVAR57<=32'b0;
	TEMP_COVAR58<=32'b0;
	TEMP_COVAR66<=32'b0;
	TEMP_COVAR67<=32'b0;
	TEMP_COVAR68<=32'b0;
	TEMP_COVAR77<=32'b0;
	TEMP_COVAR78<=32'b0;
	TEMP_COVAR88<=32'b0;




	TRIGSHIFT<=2'b0;
	DATA_READY<=0;
	COUNTER=8'b0;
end

always @(posedge M_CLK) begin
	TRIGSHIFT<={TRIGSHIFT[0],TRIGGER};
	if (TRIGSHIFT[0]&&!TRIGSHIFT[1])  begin
	   DATA_READY<=0;
		COUNTER<=8'b0;
		DATA1<=NEW_DATA1;
		DATA2<=NEW_DATA2;
		DATA3<=NEW_DATA3;
		DATA4<=NEW_DATA4;
		DATA5<=NEW_DATA5;
		DATA6<=NEW_DATA6;
		DATA7<=NEW_DATA7;
		DATA8<=NEW_DATA8;
	end //posedge du trig

	if (COUNTER<8'd16) COUNTER<=COUNTER+1;

	 if (COUNTER==8'd2) begin //converte Delta into absolute delta and sign

		if (DATA1>=MEAN1) begin DELTA_1_NEG<=1'b0;  DELTA_ABS1<=DATA1-MEAN1; end//POSITIVE 0000000000XXX
 		else begin DELTA_1_NEG<=1'b1; DELTA_ABS1<=MEAN1-DATA1; end
		if (DATA2>=MEAN2) begin DELTA_2_NEG<=1'b0;  DELTA_ABS2<=DATA2-MEAN2; end//POSITIVE 0000000000XXX
		else begin DELTA_2_NEG<=1'b1; DELTA_ABS2<=MEAN2-DATA2; end
		if (DATA3>=MEAN3) begin DELTA_3_NEG<=1'b0;  DELTA_ABS3<=DATA3-MEAN3; end//POSITIVE 0000000000XXX
		else begin DELTA_3_NEG<=1'b1; DELTA_ABS3<=MEAN3-DATA3; end
		if (DATA4>=MEAN4) begin DELTA_4_NEG<=1'b0;  DELTA_ABS4<=DATA4-MEAN4; end//POSITIVE 0000000000XXX
		else begin DELTA_4_NEG<=1'b1; DELTA_ABS4<=MEAN4-DATA4; end
		if (DATA5>=MEAN5) begin DELTA_5_NEG<=1'b0;  DELTA_ABS5<=DATA5-MEAN5; end//POSITIVE 0000000000XXX
		else begin DELTA_5_NEG<=1'b1; DELTA_ABS5<=MEAN5-DATA5; end
		if (DATA6>=MEAN6) begin DELTA_6_NEG<=1'b0;  DELTA_ABS6<=DATA6-MEAN6; end//POSITIVE 0000000000XXX
		else begin DELTA_6_NEG<=1'b1; DELTA_ABS6<=MEAN6-DATA6; end
		if (DATA7>=MEAN7) begin DELTA_7_NEG<=1'b0;  DELTA_ABS7<=DATA7-MEAN7; end//POSITIVE 0000000000XXX
		else begin DELTA_7_NEG<=1'b1; DELTA_ABS7<=MEAN7-DATA7; end
		if (DATA8>=MEAN8) begin DELTA_8_NEG<=1'b0;  DELTA_ABS8<=DATA8-MEAN8; end//POSITIVE 0000000000XXX
		else begin DELTA_8_NEG<=1'b1; DELTA_ABS8<=MEAN8-DATA8; end

	end


	else if (COUNTER==8'd3) begin //COMPUTE TEMP_MEAN  //proper way to do exponential smoothing without truncature. Always multiply positive numbers
	if (DELTA_1_NEG==0) TEMP_MEAN1<=TEMP_MEAN1+ALPHA_MEAN*DELTA_ABS1; //POSITIVE 0000000000XXX
	else TEMP_MEAN1<=TEMP_MEAN1-ALPHA_MEAN*DELTA_ABS1;//POSITIVE 0000000000XXX
	if (DELTA_2_NEG==0) TEMP_MEAN2<=TEMP_MEAN2+ALPHA_MEAN*DELTA_ABS2; //POSITIVE 0000000000XXX
	else TEMP_MEAN2<=TEMP_MEAN2-ALPHA_MEAN*DELTA_ABS2;//POSITIVE 0000000000XXX
	if (DELTA_3_NEG==0) TEMP_MEAN3<=TEMP_MEAN3+ALPHA_MEAN*DELTA_ABS3; //POSITIVE 0000000000XXX
	else TEMP_MEAN3<=TEMP_MEAN3-ALPHA_MEAN*DELTA_ABS3;//POSITIVE 0000000000XXX
	if (DELTA_4_NEG==0) TEMP_MEAN4<=TEMP_MEAN4+ALPHA_MEAN*DELTA_ABS4; //POSITIVE 0000000000XXX
	else TEMP_MEAN4<=TEMP_MEAN4-ALPHA_MEAN*DELTA_ABS4;//POSITIVE 0000000000XXX
	if (DELTA_5_NEG==0) TEMP_MEAN5<=TEMP_MEAN5+ALPHA_MEAN*DELTA_ABS5; //POSITIVE 0000000000XXX
	else TEMP_MEAN5<=TEMP_MEAN5-ALPHA_MEAN*DELTA_ABS5;//POSITIVE 0000000000XXX
	if (DELTA_6_NEG==0) TEMP_MEAN6<=TEMP_MEAN6+ALPHA_MEAN*DELTA_ABS6; //POSITIVE 0000000000XXX
	else TEMP_MEAN6<=TEMP_MEAN6-ALPHA_MEAN*DELTA_ABS6;//POSITIVE 0000000000XXX
	if (DELTA_7_NEG==0) TEMP_MEAN7<=TEMP_MEAN7+ALPHA_MEAN*DELTA_ABS7; //POSITIVE 0000000000XXX
	else TEMP_MEAN7<=TEMP_MEAN7-ALPHA_MEAN*DELTA_ABS7;//POSITIVE 0000000000XXX
	if (DELTA_8_NEG==0) TEMP_MEAN8<=TEMP_MEAN8+ALPHA_MEAN*DELTA_ABS8; //POSITIVE 0000000000XXX
	else TEMP_MEAN8<=TEMP_MEAN8-ALPHA_MEAN*DELTA_ABS8;//POSITIVE 0000000000XXX

	end

	else if (COUNTER==8'd4) begin //lets compute absolute covariance
		S11<=DELTA_ABS1*DELTA_ABS1;
		S12<=DELTA_ABS1*DELTA_ABS2;
		S13<=DELTA_ABS1*DELTA_ABS3;
		S14<=DELTA_ABS1*DELTA_ABS4;
		S15<=DELTA_ABS1*DELTA_ABS5;
		S16<=DELTA_ABS1*DELTA_ABS6;
		S17<=DELTA_ABS1*DELTA_ABS7;
		S18<=DELTA_ABS1*DELTA_ABS8;
		S22<=DELTA_ABS2*DELTA_ABS2;
		S23<=DELTA_ABS2*DELTA_ABS3;
		S24<=DELTA_ABS2*DELTA_ABS4;
		S25<=DELTA_ABS2*DELTA_ABS5;
		S26<=DELTA_ABS2*DELTA_ABS6;
		S27<=DELTA_ABS2*DELTA_ABS7;
		S28<=DELTA_ABS2*DELTA_ABS8;
		S33<=DELTA_ABS3*DELTA_ABS3;
		S34<=DELTA_ABS3*DELTA_ABS4;
		S35<=DELTA_ABS3*DELTA_ABS5;
		S36<=DELTA_ABS3*DELTA_ABS6;
		S37<=DELTA_ABS3*DELTA_ABS7;
		S38<=DELTA_ABS3*DELTA_ABS8;
		S44<=DELTA_ABS4*DELTA_ABS4;
		S45<=DELTA_ABS4*DELTA_ABS5;
		S46<=DELTA_ABS4*DELTA_ABS6;
		S47<=DELTA_ABS4*DELTA_ABS7;
		S48<=DELTA_ABS4*DELTA_ABS8;
		S55<=DELTA_ABS5*DELTA_ABS5;
		S56<=DELTA_ABS5*DELTA_ABS6;
		S57<=DELTA_ABS5*DELTA_ABS7;
		S58<=DELTA_ABS5*DELTA_ABS8;
		S66<=DELTA_ABS6*DELTA_ABS6;
		S67<=DELTA_ABS6*DELTA_ABS7;
		S68<=DELTA_ABS6*DELTA_ABS8;
		S77<=DELTA_ABS7*DELTA_ABS7;
		S78<=DELTA_ABS7*DELTA_ABS7;
		S88<=DELTA_ABS8*DELTA_ABS8;
	end

//need to reverse complement ?
//first multiply by alpha RMS ? not necessarily

	else if (COUNTER==8'd5) begin //l
		if (DELTA_1_NEG ^ DELTA_1_NEG) S11<= ~S11+1; //equivalent to -S11
		if (DELTA_1_NEG ^ DELTA_2_NEG) S12<= ~S12+1;
		if (DELTA_1_NEG ^ DELTA_3_NEG) S13<= ~S13+1;
		if (DELTA_1_NEG ^ DELTA_4_NEG) S14<= ~S14+1;
		if (DELTA_1_NEG ^ DELTA_5_NEG) S15<= ~S15+1;
		if (DELTA_1_NEG ^ DELTA_6_NEG) S16<= ~S16+1;
		if (DELTA_1_NEG ^ DELTA_7_NEG) S17<= ~S17+1;
		if (DELTA_1_NEG ^ DELTA_8_NEG) S18<= ~S18+1;

		if (DELTA_2_NEG ^ DELTA_2_NEG) S22<= ~S22+1;
		if (DELTA_2_NEG ^ DELTA_3_NEG) S23<= ~S23+1;
		if (DELTA_2_NEG ^ DELTA_4_NEG) S24<= ~S24+1;
		if (DELTA_2_NEG ^ DELTA_5_NEG) S25<= ~S25+1;
		if (DELTA_2_NEG ^ DELTA_6_NEG) S26<= ~S26+1;
		if (DELTA_2_NEG ^ DELTA_7_NEG) S27<= ~S27+1;
		if (DELTA_2_NEG ^ DELTA_8_NEG) S28<= ~S28+1;

		if (DELTA_3_NEG ^ DELTA_3_NEG) S33<= ~S33+1;
		if (DELTA_3_NEG ^ DELTA_4_NEG) S34<= ~S34+1;
		if (DELTA_3_NEG ^ DELTA_5_NEG) S35<= ~S35+1;
		if (DELTA_3_NEG ^ DELTA_6_NEG) S36<= ~S36+1;
		if (DELTA_3_NEG ^ DELTA_7_NEG) S37<= ~S37+1;
		if (DELTA_3_NEG ^ DELTA_8_NEG) S38<= ~S38+1;

		if (DELTA_4_NEG ^ DELTA_4_NEG) S44<= ~S44+1;
		if (DELTA_4_NEG ^ DELTA_5_NEG) S45<= ~S45+1;
		if (DELTA_4_NEG ^ DELTA_6_NEG) S46<= ~S46+1;
		if (DELTA_4_NEG ^ DELTA_7_NEG) S47<= ~S47+1;
		if (DELTA_4_NEG ^ DELTA_8_NEG) S48<= ~S48+1;

		if (DELTA_5_NEG ^ DELTA_5_NEG) S55<= ~S55+1;
		if (DELTA_5_NEG ^ DELTA_6_NEG) S56<= ~S56+1;
		if (DELTA_5_NEG ^ DELTA_7_NEG) S57<= ~S57+1;
		if (DELTA_5_NEG ^ DELTA_8_NEG) S58<= ~S58+1;

		if (DELTA_6_NEG ^ DELTA_6_NEG) S66<= ~S66+1;
		if (DELTA_6_NEG ^ DELTA_7_NEG) S67<= ~S67+1;
		if (DELTA_6_NEG ^ DELTA_8_NEG) S68<= ~S68+1;

		if (DELTA_7_NEG ^ DELTA_7_NEG) S77<= ~S77+1;
		if (DELTA_7_NEG ^ DELTA_8_NEG) S78<= ~S78+1;

		if (DELTA_8_NEG ^ DELTA_8_NEG) S88<= ~S88+1;

	end

	else if (COUNTER==8'd6) begin
		if (S11[15:0]>=COVAR11) TEMP_COVAR11<=TEMP_COVAR11+ALPHA_RMS*(S11[15:0]-COVAR11);
		else TEMP_COVAR11<=TEMP_COVAR11-ALPHA_RMS*(COVAR11-S11[15:0]);
	//	if (S12[15:0]>=COVAR12) TEMP_COVAR12<=TEMP_COVAR12+ALPHA_RMS*(S12[15:0]-COVAR12);
	//	else TEMP_COVAR12<=TEMP_COVAR12-ALPHA_RMS*(COVAR12-S12[15:0]);
/*		if (S13[15:0]>=COVAR13) TEMP_COVAR13<=TEMP_COVAR13+ALPHA_RMS*(S13[15:0]-COVAR13);
		else TEMP_COVAR13<=TEMP_COVAR13-ALPHA_RMS*(COVAR13-S13[15:0]);
		if (S14[15:0]>=COVAR14) TEMP_COVAR14<=TEMP_COVAR14+ALPHA_RMS*(S14[15:0]-COVAR14);
		else TEMP_COVAR14<=TEMP_COVAR14-ALPHA_RMS*(COVAR14-S14[15:0]);
		if (S15[15:0]>=COVAR15) TEMP_COVAR15<=TEMP_COVAR15+ALPHA_RMS*(S15[15:0]-COVAR15);
		else TEMP_COVAR15<=TEMP_COVAR15-ALPHA_RMS*(COVAR15-S15[15:0]);
		if (S16[15:0]>=COVAR16) TEMP_COVAR16<=TEMP_COVAR16+ALPHA_RMS*(S16[15:0]-COVAR16);
		else TEMP_COVAR16<=TEMP_COVAR16-ALPHA_RMS*(COVAR16-S16[15:0]);
		if (S17[15:0]>=COVAR17) TEMP_COVAR17<=TEMP_COVAR17+ALPHA_RMS*(S17[15:0]-COVAR17);
		else TEMP_COVAR17<=TEMP_COVAR17-ALPHA_RMS*(COVAR17-S17[15:0]);
		if (S18[15:0]>=COVAR18) TEMP_COVAR18<=TEMP_COVAR18+ALPHA_RMS*(S18[15:0]-COVAR18);
		else TEMP_COVAR18<=TEMP_COVAR18-ALPHA_RMS*(COVAR18-S18[15:0]);
*/
		if (S22[15:0]>=COVAR22) TEMP_COVAR22<=TEMP_COVAR22+ALPHA_RMS*(S22[15:0]-COVAR22);
		else TEMP_COVAR22<=TEMP_COVAR22-ALPHA_RMS*(COVAR22-S22[15:0]);
/*		if (S23[15:0]>=COVAR23) TEMP_COVAR23<=TEMP_COVAR23+ALPHA_RMS*(S23[15:0]-COVAR23);
		else TEMP_COVAR23<=TEMP_COVAR23-ALPHA_RMS*(COVAR23-S23[15:0]);
		if (S24[15:0]>=COVAR24) TEMP_COVAR24<=TEMP_COVAR24+ALPHA_RMS*(S24[15:0]-COVAR24);
		else TEMP_COVAR24<=TEMP_COVAR24-ALPHA_RMS*(COVAR24-S24[15:0]);
		if (S25[15:0]>=COVAR25) TEMP_COVAR25<=TEMP_COVAR25+ALPHA_RMS*(S25[15:0]-COVAR25);
		else TEMP_COVAR25<=TEMP_COVAR25-ALPHA_RMS*(COVAR25-S25[15:0]);
		if (S26[15:0]>=COVAR26) TEMP_COVAR26<=TEMP_COVAR26+ALPHA_RMS*(S26[15:0]-COVAR26);
		else TEMP_COVAR26<=TEMP_COVAR26-ALPHA_RMS*(COVAR26-S26[15:0]);
		if (S27[15:0]>=COVAR27) TEMP_COVAR27<=TEMP_COVAR27+ALPHA_RMS*(S27[15:0]-COVAR27);
		else TEMP_COVAR27<=TEMP_COVAR27-ALPHA_RMS*(COVAR27-S27[15:0]);
		if (S28[15:0]>=COVAR28) TEMP_COVAR28<=TEMP_COVAR28+ALPHA_RMS*(S28[15:0]-COVAR28);
		else TEMP_COVAR28<=TEMP_COVAR28-ALPHA_RMS*(COVAR28-S28[15:0]);
*/

		if (S33[15:0]>=COVAR33) TEMP_COVAR33<=TEMP_COVAR33+ALPHA_RMS*(S33[15:0]-COVAR33);
		else TEMP_COVAR33<=TEMP_COVAR33-ALPHA_RMS*(COVAR33-S33[15:0]);
/*		if (S34[15:0]>=COVAR34) TEMP_COVAR34<=TEMP_COVAR34+ALPHA_RMS*(S34[15:0]-COVAR34);
		else TEMP_COVAR34<=TEMP_COVAR34-ALPHA_RMS*(COVAR34-S34[15:0]);
		if (S35[15:0]>=COVAR35) TEMP_COVAR35<=TEMP_COVAR35+ALPHA_RMS*(S35[15:0]-COVAR35);
		else TEMP_COVAR35<=TEMP_COVAR35-ALPHA_RMS*(COVAR35-S35[15:0]);
		if (S36[15:0]>=COVAR36) TEMP_COVAR36<=TEMP_COVAR36+ALPHA_RMS*(S36[15:0]-COVAR36);
		else TEMP_COVAR36<=TEMP_COVAR36-ALPHA_RMS*(COVAR36-S36[15:0]);
		if (S37[15:0]>=COVAR37) TEMP_COVAR37<=TEMP_COVAR37+ALPHA_RMS*(S37[15:0]-COVAR37);
		else TEMP_COVAR37<=TEMP_COVAR37-ALPHA_RMS*(COVAR37-S37[15:0]);
		if (S38[15:0]>=COVAR38) TEMP_COVAR38<=TEMP_COVAR38+ALPHA_RMS*(S38[15:0]-COVAR38);
		else TEMP_COVAR38<=TEMP_COVAR38-ALPHA_RMS*(COVAR38-S38[15:0]);
*/
		if (S44[15:0]>=COVAR44) TEMP_COVAR44<=TEMP_COVAR44+ALPHA_RMS*(S44[15:0]-COVAR44);
		else TEMP_COVAR44<=TEMP_COVAR44-ALPHA_RMS*(COVAR44-S44[15:0]);
	/*	if (S45[15:0]>=COVAR45) TEMP_COVAR45<=TEMP_COVAR45+ALPHA_RMS*(S45[15:0]-COVAR45);
		else TEMP_COVAR45<=TEMP_COVAR45-ALPHA_RMS*(COVAR45-S45[15:0]);
		if (S46[15:0]>=COVAR46) TEMP_COVAR46<=TEMP_COVAR46+ALPHA_RMS*(S46[15:0]-COVAR46);
		else TEMP_COVAR46<=TEMP_COVAR46-ALPHA_RMS*(COVAR46-S46[15:0]);
		if (S47[15:0]>=COVAR47) TEMP_COVAR47<=TEMP_COVAR47+ALPHA_RMS*(S47[15:0]-COVAR47);
		else TEMP_COVAR47<=TEMP_COVAR47-ALPHA_RMS*(COVAR47-S47[15:0]);
		if (S48[15:0]>=COVAR48) TEMP_COVAR48<=TEMP_COVAR48+ALPHA_RMS*(S48[15:0]-COVAR48);
		else TEMP_COVAR48<=TEMP_COVAR48-ALPHA_RMS*(COVAR48-S48[15:0]);
*/
		if (S55[15:0]>=COVAR55) TEMP_COVAR55<=TEMP_COVAR55+ALPHA_RMS*(S55[15:0]-COVAR55);
		else TEMP_COVAR55<=TEMP_COVAR55-ALPHA_RMS*(COVAR55-S55[15:0]);
	/*	if (S56[15:0]>=COVAR56) TEMP_COVAR56<=TEMP_COVAR56+ALPHA_RMS*(S56[15:0]-COVAR56);
		else TEMP_COVAR56<=TEMP_COVAR56-ALPHA_RMS*(COVAR56-S56[15:0]);
		if (S57[15:0]>=COVAR57) TEMP_COVAR57<=TEMP_COVAR57+ALPHA_RMS*(S57[15:0]-COVAR57);
		else TEMP_COVAR57<=TEMP_COVAR57-ALPHA_RMS*(COVAR57-S57[15:0]);
		if (S58[15:0]>=COVAR58) TEMP_COVAR58<=TEMP_COVAR58+ALPHA_RMS*(S58[15:0]-COVAR58);
		else TEMP_COVAR58<=TEMP_COVAR58-ALPHA_RMS*(COVAR58-S58[15:0]);
*/
		if (S66[15:0]>=COVAR66) TEMP_COVAR66<=TEMP_COVAR66+ALPHA_RMS*(S66[15:0]-COVAR66);
		else TEMP_COVAR66<=TEMP_COVAR66-ALPHA_RMS*(COVAR66-S66[15:0]);
/*		if (S67[15:0]>=COVAR67) TEMP_COVAR67<=TEMP_COVAR67+ALPHA_RMS*(S67[15:0]-COVAR67);
		else TEMP_COVAR67<=TEMP_COVAR67-ALPHA_RMS*(COVAR67-S67[15:0]);
		if (S68[15:0]>=COVAR68) TEMP_COVAR68<=TEMP_COVAR68+ALPHA_RMS*(S68[15:0]-COVAR68);
		else TEMP_COVAR68<=TEMP_COVAR68-ALPHA_RMS*(COVAR68-S68[15:0]);
*/
		if (S77[15:0]>=COVAR77) TEMP_COVAR77<=TEMP_COVAR77+ALPHA_RMS*(S77[15:0]-COVAR77);
		else TEMP_COVAR77<=TEMP_COVAR77-ALPHA_RMS*(COVAR77-S77[15:0]);
/*		if (S78[15:0]>=COVAR78) TEMP_COVAR78<=TEMP_COVAR78+ALPHA_RMS*(S78[15:0]-COVAR78);
		else TEMP_COVAR78<=TEMP_COVAR78-ALPHA_RMS*(COVAR78-S78[15:0]);
*/
		if (S88[15:0]>=COVAR88) TEMP_COVAR88<=TEMP_COVAR88+ALPHA_RMS*(S88[15:0]-COVAR88);
		else TEMP_COVAR88<=TEMP_COVAR88-ALPHA_RMS*(COVAR88-S88[15:0]);
	end

	else if (COUNTER==8'd7) begin

		MEAN1<={TEMP_MEAN1[31],TEMP_MEAN1[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN2<={TEMP_MEAN2[31],TEMP_MEAN2[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN3<={TEMP_MEAN3[31],TEMP_MEAN3[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN4<={TEMP_MEAN4[31],TEMP_MEAN4[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN5<={TEMP_MEAN5[31],TEMP_MEAN5[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN6<={TEMP_MEAN6[31],TEMP_MEAN6[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN7<={TEMP_MEAN7[31],TEMP_MEAN7[29:15]}; //need to keep MSB in case of substraction (see above)
		MEAN8<={TEMP_MEAN8[31],TEMP_MEAN8[29:15]}; //need to keep MSB in case of substraction (see above)

		COVAR11<={TEMP_COVAR11[31],TEMP_COVAR11[29:15]};
/*	COVAR12<={TEMP_COVAR12[31],TEMP_COVAR12[29:15]};
		COVAR13<={TEMP_COVAR13[31],TEMP_COVAR13[29:15]};
		COVAR14<={TEMP_COVAR14[31],TEMP_COVAR14[29:15]};
		COVAR15<={TEMP_COVAR15[31],TEMP_COVAR15[29:15]};
		COVAR16<={TEMP_COVAR16[31],TEMP_COVAR16[29:15]};
		COVAR17<={TEMP_COVAR17[31],TEMP_COVAR17[29:15]};
		COVAR18<={TEMP_COVAR18[31],TEMP_COVAR18[29:15]};
*/
		COVAR22<={TEMP_COVAR22[31],TEMP_COVAR22[29:15]};
/*		COVAR23<={TEMP_COVAR23[31],TEMP_COVAR23[29:15]};
		COVAR24<={TEMP_COVAR24[31],TEMP_COVAR24[29:15]};
		COVAR25<={TEMP_COVAR25[31],TEMP_COVAR25[29:15]};
		COVAR26<={TEMP_COVAR26[31],TEMP_COVAR26[29:15]};
		COVAR27<={TEMP_COVAR27[31],TEMP_COVAR27[29:15]};
		COVAR28<={TEMP_COVAR28[31],TEMP_COVAR28[29:15]};*/

		COVAR33<={TEMP_COVAR33[31],TEMP_COVAR33[29:15]};
//		COVAR34<={TEMP_COVAR34[31],TEMP_COVAR34[29:15]};
//		COVAR35<={TEMP_COVAR35[31],TEMP_COVAR35[29:15]};
//		COVAR36<={TEMP_COVAR36[31],TEMP_COVAR36[29:15]};
//		COVAR37<={TEMP_COVAR37[31],TEMP_COVAR37[29:15]};
//		COVAR38<={TEMP_COVAR38[31],TEMP_COVAR38[29:15]};

		COVAR44<={TEMP_COVAR44[31],TEMP_COVAR44[29:15]};
//		COVAR45<={TEMP_COVAR45[31],TEMP_COVAR45[29:15]};
//		COVAR46<={TEMP_COVAR46[31],TEMP_COVAR46[29:15]};
//		COVAR47<={TEMP_COVAR47[31],TEMP_COVAR47[29:15]};
//		COVAR48<={TEMP_COVAR48[31],TEMP_COVAR48[29:15]};

		COVAR55<={TEMP_COVAR55[31],TEMP_COVAR55[29:15]};
//		COVAR56<={TEMP_COVAR56[31],TEMP_COVAR56[29:15]};
//		COVAR57<={TEMP_COVAR57[31],TEMP_COVAR57[29:15]};
//		COVAR58<={TEMP_COVAR58[31],TEMP_COVAR58[29:15]};

		COVAR66<={TEMP_COVAR66[31],TEMP_COVAR66[29:15]};
//		COVAR67<={TEMP_COVAR67[31],TEMP_COVAR67[29:15]};
//		COVAR68<={TEMP_COVAR68[31],TEMP_COVAR68[29:15]};

		COVAR77<={TEMP_COVAR77[31],TEMP_COVAR77[29:15]};
	//	COVAR78<={TEMP_COVAR78[31],TEMP_COVAR78[29:15]};

		COVAR88<={TEMP_COVAR88[31],TEMP_COVAR88[29:15]};

	end

	else if (COUNTER==8'd8) DATA_READY<=1;
	else if (COUNTER==8'd12) DATA_READY<=0;

end



endmodule
