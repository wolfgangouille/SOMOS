`timescale 1ns / 1ps

module RMSER_8(M_CLK,TRIGGER,NEW_DATA1,NEW_DATA2,NEW_DATA3,NEW_DATA4,NEW_DATA5,NEW_DATA6,NEW_DATA7,NEW_DATA8,RMS1,RMS2,RMS3,RMS4,RMS5,RMS6,RMS7,RMS8,DATA_READY);

input TRIGGER;
input [15:0] NEW_DATA1;
input [15:0] NEW_DATA2;
input [15:0] NEW_DATA3;
input [15:0] NEW_DATA4;
input [15:0] NEW_DATA5;
input [15:0] NEW_DATA6;
input [15:0] NEW_DATA7;
input [15:0] NEW_DATA8;
input M_CLK;
output [15:0] RMS1;
output [15:0] RMS2;
output [15:0] RMS3;
output [15:0] RMS4;
output [15:0] RMS5;
output [15:0] RMS6;
output [15:0] RMS7;
output [15:0] RMS8;
output DATA_READY;

reg [15:0] DATA1;
reg [15:0] DATA2;
reg [15:0] DATA3;
reg [15:0] DATA4;
reg [15:0] DATA5;
reg [15:0] DATA6;
reg [15:0] DATA7;
reg [15:0] DATA8;
reg [15:0] MEAN1;
reg [15:0] MEAN2;
reg [15:0] MEAN3;
reg [15:0] MEAN4;
reg [15:0] MEAN5;
reg [15:0] MEAN6;
reg [15:0] MEAN7;
reg [15:0] MEAN8;
reg [15:0] RMS1; 
reg [15:0] RMS2; 
reg [15:0] RMS3; 
reg [15:0] RMS4; 
reg [15:0] RMS5; 
reg [15:0] RMS6; 
reg [15:0] RMS7; 
reg [15:0] RMS8; 
reg [15:0] DELTA_ABS1; 
reg [15:0] DELTA_ABS2; 
reg [15:0] DELTA_ABS3; 
reg [15:0] DELTA_ABS4; 
reg [15:0] DELTA_ABS5; 
reg [15:0] DELTA_ABS6; 
reg [15:0] DELTA_ABS7; 
reg [15:0] DELTA_ABS8; 
reg [31:0] S1; 
reg [31:0] S2; 
reg [31:0] S3; 
reg [31:0] S4; 
reg [31:0] S5; 
reg [31:0] S6; 
reg [31:0] S7; 
reg [31:0] S8; 

reg [31:0] TEMP_MEAN1; 
reg [31:0] TEMP_MEAN2; 
reg [31:0] TEMP_MEAN3; 
reg [31:0] TEMP_MEAN4; 
reg [31:0] TEMP_MEAN5; 
reg [31:0] TEMP_MEAN6; 
reg [31:0] TEMP_MEAN7; 
reg [31:0] TEMP_MEAN8; 

reg [31:0] TEMP_RMS1;
reg [31:0] TEMP_RMS2;
reg [31:0] TEMP_RMS3;
reg [31:0] TEMP_RMS4;
reg [31:0] TEMP_RMS5;
reg [31:0] TEMP_RMS6;
reg [31:0] TEMP_RMS7;
reg [31:0] TEMP_RMS8;

reg [15:0] ALPHA_MEAN;
reg [15:0] ALPHA_RMS;

reg [1:0] TRIGSHIFT;
reg DATA_READY;

reg [7:0] COUNTER;

initial begin
	ALPHA_MEAN<=16'b0000000000000001;
	ALPHA_RMS<=16'b0000000000000100;	
	
	DATA1<=16'b0;
	DATA2<=16'b0;
	DATA3<=16'b0;
	DATA4<=16'b0;
	DATA5<=16'b0;
	DATA6<=16'b0;
	DATA7<=16'b0;
	DATA8<=16'b0;

	TEMP_MEAN1<=32'b10000000000000000000000000000000; 
	TEMP_MEAN2<=32'b10000000000000000000000000000000; 
	TEMP_MEAN3<=32'b10000000000000000000000000000000; 
	TEMP_MEAN4<=32'b10000000000000000000000000000000; 
	TEMP_MEAN5<=32'b10000000000000000000000000000000; 
	TEMP_MEAN6<=32'b10000000000000000000000000000000; 
	TEMP_MEAN7<=32'b10000000000000000000000000000000; 
	TEMP_MEAN8<=32'b10000000000000000000000000000000; 

	TEMP_RMS1<=32'b0; 
	TEMP_RMS2<=32'b0; 
	TEMP_RMS3<=32'b0; 
	TEMP_RMS4<=32'b0; 
	TEMP_RMS5<=32'b0; 
	TEMP_RMS6<=32'b0; 
	TEMP_RMS7<=32'b0; 
	TEMP_RMS8<=32'b0; 

	MEAN1<=16'b0000000000000000; 
	MEAN2<=16'b0000000000000000; 
	MEAN3<=16'b0000000000000000; 
	MEAN4<=16'b0000000000000000; 
	MEAN5<=16'b0000000000000000; 
	MEAN6<=16'b0000000000000000; 
	MEAN7<=16'b0000000000000000; 
	MEAN8<=16'b0000000000000000; 

	RMS1<=16'b0000000000000000; 
	RMS2<=16'b0000000000000000; 
	RMS3<=16'b0000000000000000; 
	RMS4<=16'b0000000000000000; 
	RMS5<=16'b0000000000000000; 
	RMS6<=16'b0000000000000000; 
	RMS7<=16'b0000000000000000; 
	RMS8<=16'b0000000000000000; 

	DELTA_ABS1<=16'b0;
	DELTA_ABS2<=16'b0;
	DELTA_ABS3<=16'b0;
	DELTA_ABS4<=16'b0;
	DELTA_ABS5<=16'b0;
	DELTA_ABS6<=16'b0;
	DELTA_ABS7<=16'b0;
	DELTA_ABS8<=16'b0;

	S1<=32'b0;
	S2<=32'b0;
	S3<=32'b0;
	S4<=32'b0;
	S5<=32'b0;
	S6<=32'b0;
	S7<=32'b0;
	S8<=32'b0;

	TRIGSHIFT<=2'b0;
	DATA_READY<=0;
	COUNTER=8'b0;
end

always @(posedge M_CLK) begin
	TRIGSHIFT<={TRIGSHIFT[0],TRIGGER};
	if (TRIGSHIFT[0]&&!TRIGSHIFT[1])  begin 
	   DATA_READY<=0;
		COUNTER<=8'b0; 
		DATA1<=NEW_DATA1; 
		DATA2<=NEW_DATA2; 
		DATA3<=NEW_DATA3; 
		DATA4<=NEW_DATA4; 
		DATA5<=NEW_DATA5; 
		DATA6<=NEW_DATA6; 
		DATA7<=NEW_DATA7; 
		DATA8<=NEW_DATA8; 
	end //posedge du trig
	
	if (COUNTER<8'd16) COUNTER<=COUNTER+1;

	 if (COUNTER==8'd2) begin //COMPUTE DELTA_ABS
		if (DATA1>=MEAN1) DELTA_ABS1<=DATA1-MEAN1; //POSITIVE 0000000000XXX
		else DELTA_ABS1<=MEAN1-DATA1; //POSITIVE 0000000000XXX
		if (DATA2>=MEAN2) DELTA_ABS2<=DATA2-MEAN2; //POSITIVE 0000000000XXX
		else DELTA_ABS2<=MEAN2-DATA2; //POSITIVE 0000000000XXX
		if (DATA3>=MEAN3) DELTA_ABS3<=DATA3-MEAN3; //POSITIVE 0000000000XXX
		else DELTA_ABS3<=MEAN3-DATA3; //POSITIVE 0000000000XXX		
		if (DATA4>=MEAN4) DELTA_ABS4<=DATA4-MEAN4; //POSITIVE 0000000000XXX
		else DELTA_ABS4<=MEAN4-DATA4; //POSITIVE 0000000000XXX
		if (DATA5>=MEAN5) DELTA_ABS5<=DATA5-MEAN5; //POSITIVE 0000000000XXX
		else DELTA_ABS5<=MEAN5-DATA5; //POSITIVE 0000000000XXX
		if (DATA6>=MEAN6) DELTA_ABS6<=DATA6-MEAN6; //POSITIVE 0000000000XXX
		else DELTA_ABS6<=MEAN6-DATA6; //POSITIVE 0000000000XXX
		if (DATA7>=MEAN7) DELTA_ABS7<=DATA7-MEAN7; //POSITIVE 0000000000XXX
		else DELTA_ABS7<=MEAN7-DATA7; //POSITIVE 0000000000XXX
		if (DATA8>=MEAN8) DELTA_ABS8<=DATA8-MEAN8; //POSITIVE 0000000000XXX
		else DELTA_ABS8<=MEAN8-DATA8; //POSITIVE 0000000000XXX

	end


	else if (COUNTER==8'd3) begin //COMPUTE TEMP_MEAN
		if (DATA1>=MEAN1) TEMP_MEAN1<=TEMP_MEAN1+ALPHA_MEAN*DELTA_ABS1; //POSITIVE 0000000000XXX
		else TEMP_MEAN1<=TEMP_MEAN1-ALPHA_MEAN*DELTA_ABS1;//POSITIVE 0000000000XXX
		if (DATA2>=MEAN2) TEMP_MEAN2<=TEMP_MEAN2+ALPHA_MEAN*DELTA_ABS2; //POSITIVE 0000000000XXX
		else TEMP_MEAN2<=TEMP_MEAN2-ALPHA_MEAN*DELTA_ABS2;//POSITIVE 0000000000XXX
		if (DATA3>=MEAN3) TEMP_MEAN3<=TEMP_MEAN3+ALPHA_MEAN*DELTA_ABS3; //POSITIVE 0000000000XXX
		else TEMP_MEAN3<=TEMP_MEAN3-ALPHA_MEAN*DELTA_ABS3;//POSITIVE 0000000000XXX
		if (DATA4>=MEAN4) TEMP_MEAN4<=TEMP_MEAN4+ALPHA_MEAN*DELTA_ABS4; //POSITIVE 0000000000XXX
		else TEMP_MEAN4<=TEMP_MEAN4-ALPHA_MEAN*DELTA_ABS4;//POSITIVE 0000000000XXX
		if (DATA5>=MEAN5) TEMP_MEAN5<=TEMP_MEAN5+ALPHA_MEAN*DELTA_ABS5; //POSITIVE 0000000000XXX
		else TEMP_MEAN5<=TEMP_MEAN5-ALPHA_MEAN*DELTA_ABS5;//POSITIVE 0000000000XXX
		if (DATA6>=MEAN6) TEMP_MEAN6<=TEMP_MEAN6+ALPHA_MEAN*DELTA_ABS6; //POSITIVE 0000000000XXX
		else TEMP_MEAN6<=TEMP_MEAN6-ALPHA_MEAN*DELTA_ABS6;//POSITIVE 0000000000XXX
		if (DATA7>=MEAN7) TEMP_MEAN7<=TEMP_MEAN7+ALPHA_MEAN*DELTA_ABS7; //POSITIVE 0000000000XXX
		else TEMP_MEAN7<=TEMP_MEAN7-ALPHA_MEAN*DELTA_ABS7;//POSITIVE 0000000000XXX
		if (DATA8>=MEAN8) TEMP_MEAN8<=TEMP_MEAN8+ALPHA_MEAN*DELTA_ABS8; //POSITIVE 0000000000XXX
		else TEMP_MEAN8<=TEMP_MEAN8-ALPHA_MEAN*DELTA_ABS8;//POSITIVE 0000000000XXX
	end

	else if (COUNTER==8'd4) begin 
		S1<=DELTA_ABS1*16'b000000000000001; //change square by normal
		S2<=DELTA_ABS2*16'b000000000000001; //change square by normal
		S3<=DELTA_ABS3*16'b000000000000001; //change square by normal
		S4<=DELTA_ABS4*16'b000000000000001; //change square by normal
		S5<=DELTA_ABS5*16'b000000000000001; //change square by normal
		S6<=DELTA_ABS6*16'b000000000000001; //change square by normal
		S7<=DELTA_ABS7*16'b000000000000001; //change square by normal
		S8<=DELTA_ABS8*16'b000000000000001; //change square by normal

	end
	else if (COUNTER==8'd5) begin
		if (S1[15:0]>=RMS1) TEMP_RMS1<=TEMP_RMS1+ALPHA_RMS*(S1[15:0]-RMS1);
		else TEMP_RMS1<=TEMP_RMS1-ALPHA_RMS*(RMS1-S1[15:0]);
		if (S2[15:0]>=RMS2) TEMP_RMS2<=TEMP_RMS2+ALPHA_RMS*(S2[15:0]-RMS2);
		else TEMP_RMS2<=TEMP_RMS2-ALPHA_RMS*(RMS2-S2[15:0]);
		if (S3[15:0]>=RMS3) TEMP_RMS3<=TEMP_RMS3+ALPHA_RMS*(S3[15:0]-RMS3);
		else TEMP_RMS3<=TEMP_RMS3-ALPHA_RMS*(RMS3-S3[15:0]);
		if (S4[15:0]>=RMS4) TEMP_RMS4<=TEMP_RMS4+ALPHA_RMS*(S4[15:0]-RMS4);
		else TEMP_RMS4<=TEMP_RMS4-ALPHA_RMS*(RMS4-S4[15:0]);
		if (S5[15:0]>=RMS5) TEMP_RMS5<=TEMP_RMS5+ALPHA_RMS*(S5[15:0]-RMS5);
		else TEMP_RMS5<=TEMP_RMS5-ALPHA_RMS*(RMS5-S5[15:0]);
		if (S6[15:0]>=RMS6) TEMP_RMS6<=TEMP_RMS6+ALPHA_RMS*(S6[15:0]-RMS6);
		else TEMP_RMS6<=TEMP_RMS6-ALPHA_RMS*(RMS6-S6[15:0]);
		if (S7[15:0]>=RMS7) TEMP_RMS7<=TEMP_RMS7+ALPHA_RMS*(S7[15:0]-RMS7);
		else TEMP_RMS7<=TEMP_RMS7-ALPHA_RMS*(RMS7-S7[15:0]);
		if (S8[15:0]>=RMS8) TEMP_RMS8<=TEMP_RMS8+ALPHA_RMS*(S8[15:0]-RMS8);
		else TEMP_RMS8<=TEMP_RMS8-ALPHA_RMS*(RMS8-S8[15:0]);
	end

	else if (COUNTER==8'd6) begin
		MEAN1<={TEMP_MEAN1[31],TEMP_MEAN1[29:15]}; //need to keep MSB in case of substraction (see above)
	   MEAN2<={TEMP_MEAN2[31],TEMP_MEAN2[29:15]}; 
	   MEAN3<={TEMP_MEAN3[31],TEMP_MEAN3[29:15]}; 
	   MEAN4<={TEMP_MEAN4[31],TEMP_MEAN4[29:15]}; 
	   MEAN5<={TEMP_MEAN5[31],TEMP_MEAN5[29:15]}; 
	   MEAN6<={TEMP_MEAN6[31],TEMP_MEAN6[29:15]}; 
	   MEAN7<={TEMP_MEAN7[31],TEMP_MEAN7[29:15]}; 
	   MEAN8<={TEMP_MEAN8[31],TEMP_MEAN8[29:15]}; 

		RMS1<={TEMP_RMS1[31],TEMP_RMS1[29:15]};
		RMS2<={TEMP_RMS2[31],TEMP_RMS2[29:15]};
		RMS3<={TEMP_RMS3[31],TEMP_RMS3[29:15]};
		RMS4<={TEMP_RMS4[31],TEMP_RMS4[29:15]};
		RMS5<={TEMP_RMS5[31],TEMP_RMS5[29:15]};
		RMS6<={TEMP_RMS6[31],TEMP_RMS6[29:15]};
		RMS7<={TEMP_RMS7[31],TEMP_RMS7[29:15]};
		RMS8<={TEMP_RMS8[31],TEMP_RMS8[29:15]};

	end

	else if (COUNTER==8'd7) DATA_READY<=1;
	else if (COUNTER==8'd12) DATA_READY<=0;

end



endmodule
